-------------------------------------------------------------------------------
--
-- Title       : No Title
-- Design      : Comparador4
-- Author      : Carls13
-- Company     : Carlos Hernandez
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\Admin\Desktop\Logica\Pr�cticas de Laboratorio\Pr�ctica #03\Comparador4\Comparador4\Comparador4\compile\comparador4.vhd
-- Generated   : Wed Feb 20 22:04:58 2019
-- From        : C:\Users\Admin\Desktop\Logica\Pr�cticas de Laboratorio\Pr�ctica #03\Comparador4\Comparador4\Comparador4\src\comparador4.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;

entity Comparador4 is 
end Comparador4;

architecture Comparador4 of Comparador4 is

begin

end Comparador4;
